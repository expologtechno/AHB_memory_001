`include "test.sv"
`include "idle_test.sv"
`include "mul_w_test.sv"
`include "reset_test.sv"
`include "sanity_test.sv"
`include "w_r_test.sv"
`include "wait_test.sv"
`include "size_test.sv"
`include "size0_test.sv"
`include "size1_test.sv"
`include "mem_full_test.sv"
`include "trans_test.sv"
`include "base_test.sv"
`include "arb_test.sv"
`include "error_test.sv"
`include "dummy_test.sv"
`include "w_r_constraint_test.sv"
