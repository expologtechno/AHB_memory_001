`include "sequence.sv"
`include "wait_seq.sv"
`include "idle_seq.sv"
`include "mul_wr_seq.sv"
`include "sanity_seq.sv"
`include "w_r_seq.sv"
`include "reset_seq.sv"
`include "size_seq.sv"
`include "size0_seq.sv"
`include "mem_full_seq.sv"
`include "size1_seq.sv"
`include "trans_seq.sv"
